// Code your testbench here
// or browse Examples
`timescale 1ns/1ps

//`include"testbench.v"

module tb_arithmeticologic();

	tb TB();
	
	initial begin 

		TB.pc = 32'b0;
    TB.top_CoreMem_inst.mem_instr_inst.initializeinstrMem;
    TB.iniinstrMem;
		// Initialize registers
		TB.clk = 1'b0;
		TB.rst_n = 1'b0;
		#100
		
		// Load memory
		//$readmemb("data/instrramMem_b.mem", TB.top_CoreMem_inst.mem_instr_inst.mem, 0, 3);
		$readmemh("../data/dataMem_h.mem", TB.top_CoreMem_inst.mem_data_inst.mem, 0, 3);
		
		TB.test_add;
	  TB.rst_n = 1'b0;
		#100
		
		TB.test_and;
		TB.rst_n = 1'b0;
		#100

		TB.test_andi;
		#100
    TB.rst_n = 1'b0;
    #100
		TB.test_slli;
		#100
    TB.rst_n = 1'b0;
    #100
		TB.test_slti;
		#100
    TB.rst_n = 1'b0;
    #100
		TB.test_sltiu;
  #1000
	$finish;
end

endmodule   